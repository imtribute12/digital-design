module tb();

reg [15:0] in;

wire [3:0] s_out;
wire c_out;

encoder enc(in, s_out, c_out);

initial
	begin
		in = 16'b0000_0000_0000_0001;
		#100
		in = 16'b0000_0000_0000_0010;
		#100
		in = 16'b0000_0000_0000_0100;
		#100
		in = 16'b0000_0000_0000_1000;
		#100

		in = 16'b0000_0000_0001_0000;
		#100
		in = 16'b0000_0000_0010_0000;
		#100
		in = 16'b0000_0000_0100_0000;
		#100
		in = 16'b0000_0000_1000_0000;
		#100

		in = 16'b0000_0001_0000_0000;
		#100
		in = 16'b0000_0010_0000_0000;
		#100
		in = 16'b0000_0100_0000_0000;
		#100
		in = 16'b0000_1000_0000_0000;
		#100

		in = 16'b0001_0000_0000_0000;
		#100
		in = 16'b0010_0000_0000_0000;
		#100
		in = 16'b0100_0000_0000_0000;
		#100
		in = 16'b1000_0000_0000_0000;
	end	
endmodule